`timescale 1ns/1ps

module Multiplier_4bit_t(a, b, p);

    reg [3:0] a = 4'b0;
    reg [3:0] b = 4'b0;
    wire [7:0] p;

    Multiplier_4bit(
        a.(a), 
        b.(b), 
        p.(p)
    );


    initial begin
        repeat (2 ** 4) begin
            #5 a = a + 1'b1; b = 1'b0;
            test();
            repeat (2 ** 4) begin
                #1 b = b + 1'b1;
                test();
            end
        end
        #5 $finish;
    end

    task test;
    reg [7:0] res;
    begin
        if(p != res) begin
            $display("[ERROR]");
            $write("a: %d\n", a);
            $write("b: %d\n", b);
            $write("WRONG p: %d\n", p);
            $write("SUPPOSED p: %d\n", res);
            $display;
        end
        res = a*b;
    end
    endtask

endmodule


/*
 #10 a=4'b0000; b=4'b0000;
        #10 a=4'b0001; b=4'b0000;
        #10 a=4'b0010; b=4'b0000;
        #10 a=4'b0011; b=4'b0000;
        #10 a=4'b0100; b=4'b0000;
        #10 a=4'b0101; b=4'b0000;
        #10 a=4'b0110; b=4'b0000;
        #10 a=4'b0111; b=4'b0000;
        #10 a=4'b1000; b=4'b0000;
        #10 a=4'b1001; b=4'b0000;
        #10 a=4'b1010; b=4'b0000;
        #10 a=4'b1011; b=4'b0000;
        #10 a=4'b1100; b=4'b0000;
        #10 a=4'b1101; b=4'b0000;
        #10 a=4'b1110; b=4'b0000;
        #10 a=4'b1111; b=4'b0000;

        #10 a=4'b0000; b=4'b0001;
        #10 a=4'b0001; b=4'b0001;
        #10 a=4'b0010; b=4'b0001;
        #10 a=4'b0011; b=4'b0001;
        #10 a=4'b0100; b=4'b0001;
        #10 a=4'b0101; b=4'b0001;
        #10 a=4'b0110; b=4'b0001;
        #10 a=4'b0111; b=4'b0001;
        #10 a=4'b1000; b=4'b0001;
        #10 a=4'b1001; b=4'b0001;
        #10 a=4'b1010; b=4'b0001;
        #10 a=4'b1011; b=4'b0001;
        #10 a=4'b1100; b=4'b0001;
        #10 a=4'b1101; b=4'b0001;
        #10 a=4'b1110; b=4'b0001;
        #10 a=4'b1111; b=4'b0001;

        #10 a=4'b0000; b=4'b0010;
        #10 a=4'b0001; b=4'b0010;
        #10 a=4'b0010; b=4'b0010;
        #10 a=4'b0011; b=4'b0010;
        #10 a=4'b0100; b=4'b0010;
        #10 a=4'b0101; b=4'b0010;
        #10 a=4'b0110; b=4'b0010;
        #10 a=4'b0111; b=4'b0010;
        #10 a=4'b1000; b=4'b0010;
        #10 a=4'b1001; b=4'b0010;
        #10 a=4'b1010; b=4'b0010;
        #10 a=4'b1011; b=4'b0010;
        #10 a=4'b1100; b=4'b0010;
        #10 a=4'b1101; b=4'b0010;
        #10 a=4'b1110; b=4'b0010;
        #10 a=4'b1111; b=4'b0010;

        #10 a=4'b0000; b=4'b0011;
        #10 a=4'b0001; b=4'b0011;
        #10 a=4'b0010; b=4'b0011;
        #10 a=4'b0011; b=4'b0011;
        #10 a=4'b0100; b=4'b0011;
        #10 a=4'b0101; b=4'b0011;
        #10 a=4'b0110; b=4'b0011;
        #10 a=4'b0111; b=4'b0011;
        #10 a=4'b1000; b=4'b0011;
        #10 a=4'b1001; b=4'b0011;
        #10 a=4'b1010; b=4'b0011;
        #10 a=4'b1011; b=4'b0011;
        #10 a=4'b1100; b=4'b0011;
        #10 a=4'b1101; b=4'b0011;
        #10 a=4'b1110; b=4'b0011;
        #10 a=4'b1111; b=4'b0011;

        #10 a=4'b0000; b=4'b0100;
        #10 a=4'b0001; b=4'b0100;
        #10 a=4'b0010; b=4'b0100;
        #10 a=4'b0011; b=4'b0100;
        #10 a=4'b0100; b=4'b0100;
        #10 a=4'b0101; b=4'b0100;
        #10 a=4'b0110; b=4'b0100;
        #10 a=4'b0111; b=4'b0100;
        #10 a=4'b1000; b=4'b0100;
        #10 a=4'b1001; b=4'b0100;
        #10 a=4'b1010; b=4'b0100;
        #10 a=4'b1011; b=4'b0100;
        #10 a=4'b1100; b=4'b0100;
        #10 a=4'b1101; b=4'b0100;
        #10 a=4'b1110; b=4'b0100;
        #10 a=4'b1111; b=4'b0100;

        #10 a=4'b0000; b=4'b0101;
        #10 a=4'b0001; b=4'b0101;
        #10 a=4'b0010; b=4'b0101;
        #10 a=4'b0011; b=4'b0101;
        #10 a=4'b0100; b=4'b0101;
        #10 a=4'b0101; b=4'b0101;
        #10 a=4'b0110; b=4'b0101;
        #10 a=4'b0111; b=4'b0101;
        #10 a=4'b1000; b=4'b0101;
        #10 a=4'b1001; b=4'b0101;
        #10 a=4'b1010; b=4'b0101;
        #10 a=4'b1011; b=4'b0101;
        #10 a=4'b1100; b=4'b0101;
        #10 a=4'b1101; b=4'b0101;
        #10 a=4'b1110; b=4'b0101;
        #10 a=4'b1111; b=4'b0101;

        #10 a=4'b0000; b=4'b0110;
        #10 a=4'b0001; b=4'b0110;
        #10 a=4'b0010; b=4'b0110;
        #10 a=4'b0011; b=4'b0110;
        #10 a=4'b0100; b=4'b0110;
        #10 a=4'b0101; b=4'b0110;
        #10 a=4'b0110; b=4'b0110;
        #10 a=4'b0111; b=4'b0110;
        #10 a=4'b1000; b=4'b0110;
        #10 a=4'b1001; b=4'b0110;
        #10 a=4'b1010; b=4'b0110;
        #10 a=4'b1011; b=4'b0110;
        #10 a=4'b1100; b=4'b0110;
        #10 a=4'b1101; b=4'b0110;
        #10 a=4'b1110; b=4'b0110;
        #10 a=4'b1111; b=4'b0110;

        #10 a=4'b0000; b=4'b0111;
        #10 a=4'b0001; b=4'b0111;
        #10 a=4'b0010; b=4'b0111;
        #10 a=4'b0011; b=4'b0111;
        #10 a=4'b0100; b=4'b0111;
        #10 a=4'b0101; b=4'b0111;
        #10 a=4'b0110; b=4'b0111;
        #10 a=4'b0111; b=4'b0111;
        #10 a=4'b1000; b=4'b0111;
        #10 a=4'b1001; b=4'b0111;
        #10 a=4'b1010; b=4'b0111;
        #10 a=4'b1011; b=4'b0111;
        #10 a=4'b1100; b=4'b0111;
        #10 a=4'b1101; b=4'b0111;
        #10 a=4'b1110; b=4'b0111;
        #10 a=4'b1111; b=4'b0111;
        
        #10 a=4'b0000; b=4'b1000;
        #10 a=4'b0001; b=4'b1000;
        #10 a=4'b0010; b=4'b1000;
        #10 a=4'b0011; b=4'b1000;
        #10 a=4'b0100; b=4'b1000;
        #10 a=4'b0101; b=4'b1000;
        #10 a=4'b0110; b=4'b1000;
        #10 a=4'b0111; b=4'b1000;
        #10 a=4'b1000; b=4'b1000;
        #10 a=4'b1001; b=4'b1000;
        #10 a=4'b1010; b=4'b1000;
        #10 a=4'b1011; b=4'b1000;
        #10 a=4'b1100; b=4'b1000;
        #10 a=4'b1101; b=4'b1000;
        #10 a=4'b1110; b=4'b1000;
        #10 a=4'b1111; b=4'b1000;

        #10 a=4'b0000; b=4'b1001;
        #10 a=4'b0001; b=4'b1001;
        #10 a=4'b0010; b=4'b1001;
        #10 a=4'b0011; b=4'b1001;
        #10 a=4'b0100; b=4'b1001;
        #10 a=4'b0101; b=4'b1001;
        #10 a=4'b0110; b=4'b1001;
        #10 a=4'b0111; b=4'b1001;
        #10 a=4'b1000; b=4'b1001;
        #10 a=4'b1001; b=4'b1001;
        #10 a=4'b1010; b=4'b1001;
        #10 a=4'b1011; b=4'b1001;
        #10 a=4'b1100; b=4'b1001;
        #10 a=4'b1101; b=4'b1001;
        #10 a=4'b1110; b=4'b1001;
        #10 a=4'b1111; b=4'b1001;

        #10 a=4'b0000; b=4'b1010;
        #10 a=4'b0001; b=4'b1010;
        #10 a=4'b0010; b=4'b1010;
        #10 a=4'b0011; b=4'b1010;
        #10 a=4'b0100; b=4'b1010;
        #10 a=4'b0101; b=4'b1010;
        #10 a=4'b0110; b=4'b1010;
        #10 a=4'b0111; b=4'b1010;
        #10 a=4'b1000; b=4'b1010;
        #10 a=4'b1001; b=4'b1010;
        #10 a=4'b1010; b=4'b1010;
        #10 a=4'b1011; b=4'b1010;
        #10 a=4'b1100; b=4'b1010;
        #10 a=4'b1101; b=4'b1010;
        #10 a=4'b1110; b=4'b1010;
        #10 a=4'b1111; b=4'b1010;

        #10 a=4'b0000; b=4'b1011;
        #10 a=4'b0001; b=4'b1011;
        #10 a=4'b0010; b=4'b1011;
        #10 a=4'b0011; b=4'b1011;
        #10 a=4'b0100; b=4'b1011;
        #10 a=4'b0101; b=4'b1011;
        #10 a=4'b0110; b=4'b1011;
        #10 a=4'b0111; b=4'b1011;
        #10 a=4'b1000; b=4'b1011;
        #10 a=4'b1001; b=4'b1011;
        #10 a=4'b1010; b=4'b1011;
        #10 a=4'b1011; b=4'b1011;
        #10 a=4'b1100; b=4'b1011;
        #10 a=4'b1101; b=4'b1011;
        #10 a=4'b1110; b=4'b1011;
        #10 a=4'b1111; b=4'b1011;

        #10 a=4'b0000; b=4'b1100;
        #10 a=4'b0001; b=4'b1100;
        #10 a=4'b0010; b=4'b1100;
        #10 a=4'b0011; b=4'b1100;
        #10 a=4'b0100; b=4'b1100;
        #10 a=4'b0101; b=4'b1100;
        #10 a=4'b0110; b=4'b1100;
        #10 a=4'b0111; b=4'b1100;
        #10 a=4'b1000; b=4'b1100;
        #10 a=4'b1001; b=4'b1100;
        #10 a=4'b1010; b=4'b1100;
        #10 a=4'b1011; b=4'b1100;
        #10 a=4'b1100; b=4'b1100;
        #10 a=4'b1101; b=4'b1100;
        #10 a=4'b1110; b=4'b1100;
        #10 a=4'b1111; b=4'b1100;

        #10 a=4'b0000; b=4'b1101;
        #10 a=4'b0001; b=4'b1101;
        #10 a=4'b0010; b=4'b1101;
        #10 a=4'b0011; b=4'b1101;
        #10 a=4'b0100; b=4'b1101;
        #10 a=4'b0101; b=4'b1101;
        #10 a=4'b0110; b=4'b1101;
        #10 a=4'b0111; b=4'b1101;
        #10 a=4'b1000; b=4'b1101;
        #10 a=4'b1001; b=4'b1101;
        #10 a=4'b1010; b=4'b1101;
        #10 a=4'b1011; b=4'b1101;
        #10 a=4'b1100; b=4'b1101;
        #10 a=4'b1101; b=4'b1101;
        #10 a=4'b1110; b=4'b1101;
        #10 a=4'b1111; b=4'b1101;

        #10 a=4'b0000; b=4'b1110;
        #10 a=4'b0001; b=4'b1110;
        #10 a=4'b0010; b=4'b1110;
        #10 a=4'b0011; b=4'b1110;
        #10 a=4'b0100; b=4'b1110;
        #10 a=4'b0101; b=4'b1110;
        #10 a=4'b0110; b=4'b1110;
        #10 a=4'b0111; b=4'b1110;
        #10 a=4'b1000; b=4'b1110;
        #10 a=4'b1001; b=4'b1110;
        #10 a=4'b1010; b=4'b1110;
        #10 a=4'b1011; b=4'b1110;
        #10 a=4'b1100; b=4'b1110;
        #10 a=4'b1101; b=4'b1110;
        #10 a=4'b1110; b=4'b1110;
        #10 a=4'b1111; b=4'b1110;

        #10 a=4'b0000; b=4'b1111;
        #10 a=4'b0001; b=4'b1111;
        #10 a=4'b0010; b=4'b1111;
        #10 a=4'b0011; b=4'b1111;
        #10 a=4'b0100; b=4'b1111;
        #10 a=4'b0101; b=4'b1111;
        #10 a=4'b0110; b=4'b1111;
        #10 a=4'b0111; b=4'b1111;
        #10 a=4'b1000; b=4'b1111;
        #10 a=4'b1001; b=4'b1111;
        #10 a=4'b1010; b=4'b1111;
        #10 a=4'b1011; b=4'b1111;
        #10 a=4'b1100; b=4'b1111;
        #10 a=4'b1101; b=4'b1111;
        #10 a=4'b1110; b=4'b1111;
        #10 a=4'b1111; b=4'b1111;
/*